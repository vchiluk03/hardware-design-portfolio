# Source Code Withheld

This file is intentionally withheld to comply with academic integrity and responsible sharing practices.

Project context, reports, and documentation remain available in this public repository.

Access request link: https://github.com/vchiluk03/hardware-design-portfolio/issues/new?template=code_access_request.yml&title=Code%20Access%20Request

Original path: I2CMB-Controller-Verification\project_benches\rtl\bus_state.vhd


