﻿# Source Code Withheld

This file is intentionally withheld to comply with academic integrity and responsible sharing practices.

Project context, reports, and documentation remain available in this public repository.

Access request link: https://github.com/<your-username>/<private-code-repo>/issues/new?title=Project%20Code%20Access%20Request

Original path: LC3-CPU-Decode-UVM\decode_unit_uvm\tb\tests\src\test_top.svh


